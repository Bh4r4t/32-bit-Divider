`timescale 1ns / 1ps

module comparator(
    input [31:0] a,
    input [31:0] b,
    output a_l
    );
    
    wire [31:0] E, A;
    Compare1 cp0(a[0], b[0], E[0], A[0]);
    Compare1 cp1(a[1], b[1], E[1], A[1]);
    Compare1 cp2(a[2], b[2], E[2], A[2]);
    Compare1 cp3(a[3], b[3], E[3], A[3]);
    Compare1 cp4(a[4], b[4], E[4], A[4]);
    Compare1 cp5(a[5], b[5], E[5], A[5]);
    Compare1 cp6(a[6], b[6], E[6], A[6]);
    Compare1 cp7(a[7], b[7], E[7], A[7]);
    Compare1 cp8(a[8], b[8], E[8], A[8]);
    Compare1 cp9(a[9], b[9], E[9], A[9]);
    Compare1 cp10(a[10], b[10], E[10], A[10]);
    Compare1 cp11(a[11], b[11], E[11], A[11]);
    Compare1 cp12(a[12], b[12], E[12], A[12]);
    Compare1 cp13(a[13], b[13], E[13], A[13]);
    Compare1 cp14(a[14], b[14], E[14], A[14]);
    Compare1 cp15(a[15], b[15], E[15], A[15]);
    Compare1 cp16(a[16], b[16], E[16], A[16]);
    Compare1 cp17(a[17], b[17], E[17], A[17]);
    Compare1 cp18(a[18], b[18], E[18], A[18]);
    Compare1 cp19(a[19], b[19], E[19], A[19]);
    Compare1 cp20(a[20], b[20], E[20], A[20]);
    Compare1 cp21(a[21], b[21], E[21], A[21]);
    Compare1 cp22(a[22], b[22], E[22], A[22]);
    Compare1 cp23(a[23], b[23], E[23], A[23]);
    Compare1 cp24(a[24], b[24], E[24], A[24]);
    Compare1 cp25(a[25], b[25], E[25], A[25]);
    Compare1 cp26(a[26], b[26], E[26], A[26]);
    Compare1 cp27(a[27], b[27], E[27], A[27]);
    Compare1 cp28(a[28], b[28], E[28], A[28]);
    Compare1 cp29(a[29], b[29], E[29], A[29]);
    Compare1 cp30(a[30], b[30], E[30], A[30]);
    Compare1 cp31(a[31], b[31], E[31], A[31]);
    
    
    assign a_l =  ( A[31] |
                   (A[30]&E[31]) |
                   (A[29]&E[30]&E[31]) | 
                   (A[28]&E[31]&E[30]&E[29]) |
                   (A[27]&E[31]&E[30]&E[29]&E[28]) |
                   (A[26]&E[31]&E[30]&E[29]&E[28]&E[27]) |
                   (A[25]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]) |
                   (A[24]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]) |
                   (A[23]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]) |
                   (A[22]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]) |
                   (A[21]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]) |
                   (A[20]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]) |
                   (A[19]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]) | 
                   (A[18]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]) |
                   (A[17]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]) |
                   (A[16]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]) |
                   (A[15]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]) | 
                   (A[14]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]) |
                   (A[13]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]) |
                   (A[12]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]) | 
                   (A[11]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]) |
                   (A[10]&E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]) |
                   (A[9] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]) |
                   (A[8] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]) |
                   (A[7] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]) |
                   (A[6] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]) |
                   (A[5] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]&E[6]) |
                   (A[4] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]&E[6]&E[5]) |
                   (A[3] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]&E[6]&E[5]&E[4]) |
                   (A[2] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]&E[6]&E[5]&E[4]&E[3]) |
                   (A[1] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]&E[6]&E[5]&E[4]&E[3]&E[2]) |
                   (A[0] &E[31]&E[30]&E[29]&E[28]&E[27]&E[26]&E[25]&E[24]&E[23]&E[22]&E[21]&E[20]&E[19]&E[18]&E[17]&E[16]&E[15]&E[14]&E[13]&E[12]&E[11]&E[10]&E[9]&E[8]&E[7]&E[6]&E[5]&E[4]&E[3]&E[2]&E[1])
                    );    
    
endmodule


module Compare1(
    input a,
    input b,
    output equal, 
    output a_less
    );
    
    assign equal = (a&b) | (~a & ~b);
    assign a_less = (~a & b);
        
endmodule